module mux50_1(
input clk,
input [15:0] a_1,
input [15:0] a_2,
input [15:0] a_3,
input [15:0] a_4,
input [15:0] a_5,
input [15:0] a_6,
input [15:0] a_7,
input [15:0] a_8,
input [15:0] a_9,
input [15:0] a_10,
input [15:0] a_11,
input [15:0] a_12,
input [15:0] a_13,
input [15:0] a_14,
input [15:0] a_15,
input [15:0] a_16,
input [15:0] a_17,
input [15:0] a_18,
input [15:0] a_19,
input [15:0] a_20,
input [15:0] a_21,
input [15:0] a_22,
input [15:0] a_23,
input [15:0] a_24,
input [15:0] a_25,
input [15:0] a_26,
input [15:0] a_27,
input [15:0] a_28,
input [15:0] a_29,
input [15:0] a_30,
input [15:0] a_31,
input [15:0] a_32,
input [15:0] a_33,
input [15:0] a_34,
input [15:0] a_35,
input [15:0] a_36,
input [15:0] a_37,
input [15:0] a_38,
input [15:0] a_39,
input [15:0] a_40,
input [15:0] a_41,
input [15:0] a_42,
input [15:0] a_43,
input [15:0] a_44,
input [15:0] a_45,
input [15:0] a_46,
input [15:0] a_47,
input [15:0] a_48,
input [15:0] a_49,
input [15:0] a_50,
input [15:0] a_51,
input [15:0] a_52,
input [15:0] a_53,
input [15:0] a_54,
input [15:0] a_55,
input [15:0] a_56,
input [15:0] a_57,
input [15:0] a_58,
input [15:0] a_59,
input [15:0] a_60,
input [15:0] a_61,
input [15:0] a_62,
input [15:0] a_63,
input [15:0] a_64,
input [15:0] a_65,
input [15:0] a_66,
input [15:0] a_67,
input [15:0] a_68,
input [15:0] a_69,
input [15:0] a_70,
input [15:0] a_71,
input [15:0] a_72,
input [15:0] a_73,
input [15:0] a_74,
input [15:0] a_75,
input [15:0] a_76,
input [15:0] a_77,
input [15:0] a_78,
input [15:0] a_79,
input [15:0] a_80,
input [15:0] a_81,
input [15:0] a_82,
input [15:0] a_83,
input [15:0] a_84,
input [15:0] a_85,
input [15:0] a_86,
input [15:0] a_87,
input [15:0] a_88,
input [15:0] a_89,
input [15:0] a_90,
input [15:0] a_91,
input [15:0] a_92,
input [15:0] a_93,
input [15:0] a_94,
input [15:0] a_95,
input [15:0] a_96,
input [15:0] a_97,
input [15:0] a_98,
input [15:0] a_99,
input [15:0] a_100,
input [15:0] a_101,
input [15:0] a_102,
input [15:0] a_103,
input [15:0] a_104,
input [15:0] a_105,
input [15:0] a_106,
input [15:0] a_107,
input [15:0] a_108,
input [15:0] a_109,
input [15:0] a_110,
input [15:0] a_111,
input [15:0] a_112,
input [15:0] a_113,
input [15:0] a_114,
input [15:0] a_115,
input [15:0] a_116,
input [15:0] a_117,
input [15:0] a_118,
input [15:0] a_119,
input [15:0] a_120,
input [15:0] a_121,
input [15:0] a_122,
input [15:0] a_123,
input [15:0] a_124,
input [15:0] a_125,
input [15:0] a_126,
input [15:0] a_127,
input [15:0] a_128,
input [15:0] a_129,
input [15:0] a_130,
input [15:0] a_131,
input [15:0] a_132,
input [15:0] a_133,
input [15:0] a_134,
input [15:0] a_135,
input [15:0] a_136,
input [15:0] a_137,
input [15:0] a_138,
input [15:0] a_139,
input [15:0] a_140,
input [15:0] a_141,
input [15:0] a_142,
input [15:0] a_143,
input [15:0] a_144,
input [15:0] a_145,
input [15:0] a_146,
input [15:0] a_147,
input [15:0] a_148,
input [15:0] a_149,
input [15:0] a_150,
input [15:0] a_151,
input [15:0] a_152,
input [15:0] a_153,
input [15:0] a_154,
input [15:0] a_155,
input [15:0] a_156,
input [15:0] a_157,
input [15:0] a_158,
input [15:0] a_159,
input [15:0] a_160,
input [15:0] a_161,
input [15:0] a_162,
input [15:0] a_163,
input [15:0] a_164,
input [15:0] a_165,
input [15:0] a_166,
input [15:0] a_167,
input [15:0] a_168,
input [15:0] a_169,
input [15:0] a_170,
input [15:0] a_171,
input [15:0] a_172,
input [15:0] a_173,
input [15:0] a_174,
input [15:0] a_175,
input [15:0] a_176,
input [15:0] a_177,
input [15:0] a_178,
input [15:0] a_179,
input [15:0] a_180,
input [15:0] a_181,
input [15:0] a_182,
input [15:0] a_183,
input [15:0] a_184,
input [15:0] a_185,
input [15:0] a_186,
input [15:0] a_187,
input [15:0] a_188,
input [15:0] a_189,
input [15:0] a_190,
input [15:0] a_191,
input [15:0] a_192,
input [15:0] a_193,
input [15:0] a_194,
input [15:0] a_195,
input [15:0] a_196,
input [15:0] a_197,
input [15:0] a_198,
input [15:0] a_199,
input [15:0] a_200,
input [15:0] a_201,
input [15:0] a_202,
input [15:0] a_203,
input [15:0] a_204,
input [15:0] a_205,
input [15:0] a_206,
input [15:0] a_207,
input [15:0] a_208,
input [15:0] a_209,
input [15:0] a_210,
input [15:0] a_211,
input [15:0] a_212,
input [15:0] a_213,
input [15:0] a_214,
input [15:0] a_215,
input [15:0] a_216,
input [15:0] a_217,
input [15:0] a_218,
input [15:0] a_219,
input [15:0] a_220,
input [15:0] a_221,
input [15:0] a_222,
input [15:0] a_223,
input [15:0] a_224,
input [15:0] a_225,
input [15:0] a_226,
input [15:0] a_227,
input [15:0] a_228,
input [15:0] a_229,
input [15:0] a_230,
input [15:0] a_231,
input [15:0] a_232,
input [15:0] a_233,
input [15:0] a_234,
input [15:0] a_235,
input [15:0] a_236,
input [15:0] a_237,
input [15:0] a_238,
input [15:0] a_239,
input [15:0] a_240,
input [15:0] a_241,
input [15:0] a_242,
input [15:0] a_243,
input [15:0] a_244,
input [15:0] a_245,
input [15:0] a_246,
input [15:0] a_247,
input [15:0] a_248,
input [15:0] a_249,
input [15:0] a_250,
input [15:0] a_251,
input [15:0] a_252,
input [15:0] a_253,
input [15:0] a_254,
input [15:0] a_255,
input [15:0] a_256,
input [15:0] a_257,
input [15:0] a_258,
input [15:0] a_259,
input [15:0] a_260,
input [15:0] a_261,
input [15:0] a_262,
input [15:0] a_263,
input [15:0] a_264,
input [15:0] a_265,
input [15:0] a_266,
input [15:0] a_267,
input [15:0] a_268,
input [15:0] a_269,
input [15:0] a_270,
input [15:0] a_271,
input [15:0] a_272,
input [15:0] a_273,
input [15:0] a_274,
input [15:0] a_275,
input [15:0] a_276,
input [15:0] a_277,
input [15:0] a_278,
input [15:0] a_279,
input [15:0] a_280,
input [15:0] a_281,
input [15:0] a_282,
input [15:0] a_283,
input [15:0] a_284,
input [15:0] a_285,
input [15:0] a_286,
input [15:0] a_287,
input [15:0] a_288,
output reg [15:0] ans);

reg [8:0] counter=0;
always @(posedge clk)
begin
    case (counter)
    9'h00: ans <= a_1;
    9'h01: ans <= a_2;
    9'h02: ans <= a_3;
    9'h03: ans <= a_4;
    9'h04: ans <= a_5;
    9'h05: ans <= a_6;
    9'h06: ans <= a_7;
    9'h07: ans <= a_8;
    9'h08: ans <= a_9;
    9'h09: ans <= a_10;
    9'h0A: ans <= a_11;
    9'h0B: ans <= a_12;
    9'h0C: ans <= a_13;
    9'h0D: ans <= a_14;
    9'h0E: ans <= a_15;
    9'h0F: ans <= a_16;
    9'h10: ans <= a_17;
    9'h11: ans <= a_18;
    9'h12: ans <= a_19;
    9'h13: ans <= a_20;
    9'h14: ans <= a_21;
    9'h15: ans <= a_22;
    9'h16: ans <= a_23;
    9'h17: ans <= a_24;
    9'h18: ans <= a_25;
    9'h19: ans <= a_26;
    9'h1A: ans <= a_27;
    9'h1B: ans <= a_28;
    9'h1C: ans <= a_29;
    9'h1D: ans <= a_30;
    9'h1E: ans <= a_31;
    9'h1F: ans <= a_32;
    9'h20: ans <= a_33;
    9'h21: ans <= a_34;
    9'h22: ans <= a_35;
    9'h23: ans <= a_36;
    9'h24: ans <= a_37;
    9'h25: ans <= a_38;
    9'h26: ans <= a_39;
    9'h27: ans <= a_40;
    9'h28: ans <= a_41;
    9'h29: ans <= a_42;
    9'h2A: ans <= a_43;
    9'h2B: ans <= a_44;
    9'h2C: ans <= a_45;
    9'h2D: ans <= a_46;
    9'h2E: ans <= a_47;
    9'h2F: ans <= a_48;
    9'h30: ans <= a_49;
    9'h31: ans <= a_50;
    9'h32: ans <= a_51;
    9'h33: ans <= a_52;
    9'h34: ans <= a_53;
    9'h35: ans <= a_54;
    9'h36: ans <= a_55;
    9'h37: ans <= a_56;
    9'h38: ans <= a_57;
    9'h39: ans <= a_58;
    9'h3A: ans <= a_59;
    9'h3B: ans <= a_60;
    9'h3C: ans <= a_61;
    9'h3D: ans <= a_62;
    9'h3E: ans <= a_63;
    9'h3F: ans <= a_64;
    9'h40: ans <= a_65;
    9'h41: ans <= a_66;
    9'h42: ans <= a_67;
    9'h43: ans <= a_68;
    9'h44: ans <= a_69;
    9'h45: ans <= a_70;
    9'h46: ans <= a_71;
    9'h47: ans <= a_72;
    9'h48: ans <= a_73;
    9'h49: ans <= a_74;
    9'h4A: ans <= a_75;
    9'h4B: ans <= a_76;
    9'h4C: ans <= a_77;
    9'h4D: ans <= a_78;
    9'h4E: ans <= a_79;
    9'h4F: ans <= a_80;
    9'h50: ans <= a_81;
    9'h51: ans <= a_82;
    9'h52: ans <= a_83;
    9'h53: ans <= a_84;
    9'h54: ans <= a_85;
    9'h55: ans <= a_86;
    9'h56: ans <= a_87;
    9'h57: ans <= a_88;
    9'h58: ans <= a_89;
    9'h59: ans <= a_90;
    9'h5A: ans <= a_91;
    9'h5B: ans <= a_92;
    9'h5C: ans <= a_93;
    9'h5D: ans <= a_94;
    9'h5E: ans <= a_95;
    9'h5F: ans <= a_96;
    9'h60: ans <= a_97;
    9'h61: ans <= a_98;
    9'h62: ans <= a_99;
    9'h63: ans <= a_100;
    9'h64: ans <= a_101;
    9'h65: ans <= a_102;
    9'h66: ans <= a_103;
    9'h67: ans <= a_104;
    9'h68: ans <= a_105;
    9'h69: ans <= a_106;
    9'h6A: ans <= a_107;
    9'h6B: ans <= a_108;
    9'h6C: ans <= a_109;
    9'h6D: ans <= a_110;
    9'h6E: ans <= a_111;
    9'h6F: ans <= a_112;
    9'h70: ans <= a_113;
    9'h71: ans <= a_114;
    9'h72: ans <= a_115;
    9'h73: ans <= a_116;
    9'h74: ans <= a_117;
    9'h75: ans <= a_118;
    9'h76: ans <= a_119;
    9'h77: ans <= a_120;
    9'h78: ans <= a_121;
    9'h79: ans <= a_122;
    9'h7A: ans <= a_123;
    9'h7B: ans <= a_124;
    9'h7C: ans <= a_125;
    9'h7D: ans <= a_126;
    9'h7E: ans <= a_127;
    9'h7F: ans <= a_128;
    9'h80: ans <= a_129;
    9'h81: ans <= a_130;
    9'h82: ans <= a_131;
    9'h83: ans <= a_132;
    9'h84: ans <= a_133;
    9'h85: ans <= a_134;
    9'h86: ans <= a_135;
    9'h87: ans <= a_136;
    9'h88: ans <= a_137;
    9'h89: ans <= a_138;
    9'h8A: ans <= a_139;
    9'h8B: ans <= a_140;
    9'h8C: ans <= a_141;
    9'h8D: ans <= a_142;
    9'h8E: ans <= a_143;
    9'h8F: ans <= a_144;
    9'h90: ans <= a_145;
    9'h91: ans <= a_146;
    9'h92: ans <= a_147;
    9'h93: ans <= a_148;
    9'h94: ans <= a_149;
    9'h95: ans <= a_150;
    9'h96: ans <= a_151;
    9'h97: ans <= a_152;
    9'h98: ans <= a_153;
    9'h99: ans <= a_154;
    9'h9A: ans <= a_155;
    9'h9B: ans <= a_156;
    9'h9C: ans <= a_157;
    9'h9D: ans <= a_158;
    9'h9E: ans <= a_159;
    9'h9F: ans <= a_160;
    9'hA0: ans <= a_161;
    9'hA1: ans <= a_162;
    9'hA2: ans <= a_163;
    9'hA3: ans <= a_164;
    9'hA4: ans <= a_165;
    9'hA5: ans <= a_166;
    9'hA6: ans <= a_167;
    9'hA7: ans <= a_168;
    9'hA8: ans <= a_169;
    9'hA9: ans <= a_170;
    9'hAA: ans <= a_171;
    9'hAB: ans <= a_172;
    9'hAC: ans <= a_173;
    9'hAD: ans <= a_174;
    9'hAE: ans <= a_175;
    9'hAF: ans <= a_176;
    9'hB0: ans <= a_177;
    9'hB1: ans <= a_178;
    9'hB2: ans <= a_179;
    9'hB3: ans <= a_180;
    9'hB4: ans <= a_181;
    9'hB5: ans <= a_182;
    9'hB6: ans <= a_183;
    9'hB7: ans <= a_184;
    9'hB8: ans <= a_185;
    9'hB9: ans <= a_186;
    9'hBA: ans <= a_187;
    9'hBB: ans <= a_188;
    9'hBC: ans <= a_189;
    9'hBD: ans <= a_190;
    9'hBE: ans <= a_191;
    9'hBF: ans <= a_192;
    9'hC0: ans <= a_193;
    9'hC1: ans <= a_194;
    9'hC2: ans <= a_195;
    9'hC3: ans <= a_196;
    9'hC4: ans <= a_197;
    9'hC5: ans <= a_198;
    9'hC6: ans <= a_199;
    9'hC7: ans <= a_200;
    9'hC8: ans <= a_201;
    9'hC9: ans <= a_202;
    9'hCA: ans <= a_203;
    9'hCB: ans <= a_204;
    9'hCC: ans <= a_205;
    9'hCD: ans <= a_206;
    9'hCE: ans <= a_207;
    9'hCF: ans <= a_208;
    9'hD0: ans <= a_209;
    9'hD1: ans <= a_210;
    9'hD2: ans <= a_211;
    9'hD3: ans <= a_212;
    9'hD4: ans <= a_213;
    9'hD5: ans <= a_214;
    9'hD6: ans <= a_215;
    9'hD7: ans <= a_216;
    9'hD8: ans <= a_217;
    9'hD9: ans <= a_218;
    9'hDA: ans <= a_219;
    9'hDB: ans <= a_220;
    9'hDC: ans <= a_221;
    9'hDD: ans <= a_222;
    9'hDE: ans <= a_223;
    9'hDF: ans <= a_224;
    9'hE0: ans <= a_225;
    9'hE1: ans <= a_226;
    9'hE2: ans <= a_227;
    9'hE3: ans <= a_228;
    9'hE4: ans <= a_229;
    9'hE5: ans <= a_230;
    9'hE6: ans <= a_231;
    9'hE7: ans <= a_232;
    9'hE8: ans <= a_233;
    9'hE9: ans <= a_234;
    9'hEA: ans <= a_235;
    9'hEB: ans <= a_236;
    9'hEC: ans <= a_237;
    9'hED: ans <= a_238;
    9'hEE: ans <= a_239;
    9'hEF: ans <= a_240;
    9'hF0: ans <= a_241;
    9'hF1: ans <= a_242;
    9'hF2: ans <= a_243;
    9'hF3: ans <= a_244;
    9'hF4: ans <= a_245;
    9'hF5: ans <= a_246;
    9'hF6: ans <= a_247;
    9'hF7: ans <= a_248;
    9'hF8: ans <= a_249;
    9'hF9: ans <= a_250;
    9'hFA: ans <= a_251;
    9'hFB: ans <= a_252;
    9'hFC: ans <= a_253;
    9'hFD: ans <= a_254;
    9'hFE: ans <= a_255;
    9'hFF: ans <= a_256;
    9'h100: ans <= a_257;
    9'h101: ans <= a_258;
    9'h102: ans <= a_259;
    9'h103: ans <= a_260;
    9'h104: ans <= a_261;
    9'h105: ans <= a_262;
    9'h106: ans <= a_263;
    9'h107: ans <= a_264;
    9'h108: ans <= a_265;
    9'h109: ans <= a_266;
    9'h10A: ans <= a_267;
    9'h10B: ans <= a_268;
    9'h10C: ans <= a_269;
    9'h10D: ans <= a_270;
    9'h10E: ans <= a_271;
    9'h10F: ans <= a_272;
    9'h110: ans <= a_273;
    9'h111: ans <= a_274;
    9'h112: ans <= a_275;
    9'h113: ans <= a_276;
    9'h114: ans <= a_277;
    9'h115: ans <= a_278;
    9'h116: ans <= a_279;
    9'h117: ans <= a_280;
    9'h118: ans <= a_281;
    9'h119: ans <= a_282;
    9'h11A: ans <= a_283;
    9'h11B: ans <= a_284;
    9'h11C: ans <= a_285;
    9'h11D: ans <= a_286;
    9'h11E: ans <= a_287;
    9'h11F: ans <= a_288;
    default: ans <= 9'h0; // Default value, if needed


endcase 
counter<=counter+1;
end

endmodule

