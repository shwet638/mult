module demux(input [7:0] a,
input clk,
output reg [7:0] a_1,
output reg [7:0] a_2,
output reg [7:0] a_3,
output reg [7:0] a_4,
output reg [7:0] a_5,
output reg [7:0] a_6,
output reg [7:0] a_7,
output reg [7:0] a_8,
output reg [7:0] a_9,
output reg [7:0] a_10,
output reg [7:0] a_11,
output reg [7:0] a_12,
output reg [7:0] a_13,
output reg [7:0] a_14,
output reg [7:0] a_15,
output reg [7:0] a_16,
output reg [7:0] a_17,
output reg [7:0] a_18,
output reg [7:0] a_19,
output reg [7:0] a_20,
output reg [7:0] a_21,
output reg [7:0] a_22,
output reg [7:0] a_23,
output reg [7:0] a_24,
output reg [7:0] a_25,
output reg [7:0] a_26,
output reg [7:0] a_27,
output reg [7:0] a_28,
output reg [7:0] a_29,
output reg [7:0] a_30,
output reg [7:0] a_31,
output reg [7:0] a_32,
output reg [7:0] a_33,
output reg [7:0] a_34,
output reg [7:0] a_35,
output reg [7:0] a_36,
output reg [7:0] a_37,
output reg [7:0] a_38,
output reg [7:0] a_39,
output reg [7:0] a_40,
output reg [7:0] a_41,
output reg [7:0] a_42,
output reg [7:0] a_43,
output reg [7:0] a_44,
output reg [7:0] a_45,
output reg [7:0] a_46,
output reg [7:0] a_47,
output reg [7:0] a_48,
output reg [7:0] a_49,
output reg [7:0] a_50,
output reg [7:0] a_51,
output reg [7:0] a_52,
output reg [7:0] a_53,
output reg [7:0] a_54,
output reg [7:0] a_55,
output reg [7:0] a_56,
output reg [7:0] a_57,
output reg [7:0] a_58,
output reg [7:0] a_59,
output reg [7:0] a_60,
output reg [7:0] a_61,
output reg [7:0] a_62,
output reg [7:0] a_63,
output reg [7:0] a_64,
output reg [7:0] a_65,
output reg [7:0] a_66,
output reg [7:0] a_67,
output reg [7:0] a_68,
output reg [7:0] a_69,
output reg [7:0] a_70,
output reg [7:0] a_71,
output reg [7:0] a_72,
output reg [7:0] a_73,
output reg [7:0] a_74,
output reg [7:0] a_75,
output reg [7:0] a_76,
output reg [7:0] a_77,
output reg [7:0] a_78,
output reg [7:0] a_79,
output reg [7:0] a_80,
output reg [7:0] a_81,
output reg [7:0] a_82,
output reg [7:0] a_83,
output reg [7:0] a_84,
output reg [7:0] a_85,
output reg [7:0] a_86,
output reg [7:0] a_87,
output reg [7:0] a_88,
output reg [7:0] a_89,
output reg [7:0] a_90,
output reg [7:0] a_91,
output reg [7:0] a_92,
output reg [7:0] a_93,
output reg [7:0] a_94,
output reg [7:0] a_95,
output reg [7:0] a_96,
output reg [7:0] a_97,
output reg [7:0] a_98,
output reg [7:0] a_99,
output reg [7:0] a_100,
output reg [7:0] a_101,
output reg [7:0] a_102,
output reg [7:0] a_103,
output reg [7:0] a_104,
output reg [7:0] a_105,
output reg [7:0] a_106,
output reg [7:0] a_107,
output reg [7:0] a_108,
output reg [7:0] a_109,
output reg [7:0] a_110,
output reg [7:0] a_111,
output reg [7:0] a_112,
output reg [7:0] a_113,
output reg [7:0] a_114,
output reg [7:0] a_115,
output reg [7:0] a_116,
output reg [7:0] a_117,
output reg [7:0] a_118,
output reg [7:0] a_119,
output reg [7:0] a_120,
output reg [7:0] a_121,
output reg [7:0] a_122,
output reg [7:0] a_123,
output reg [7:0] a_124,
output reg [7:0] a_125,
output reg [7:0] a_126,
output reg [7:0] a_127,
output reg [7:0] a_128,
output reg [7:0] a_129,
output reg [7:0] a_130,
output reg [7:0] a_131,
output reg [7:0] a_132,
output reg [7:0] a_133,
output reg [7:0] a_134,
output reg [7:0] a_135,
output reg [7:0] a_136,
output reg [7:0] a_137,
output reg [7:0] a_138,
output reg [7:0] a_139,
output reg [7:0] a_140,
output reg [7:0] a_141,
output reg [7:0] a_142,
output reg [7:0] a_143,
output reg [7:0] a_144,
output reg [7:0] a_145,
output reg [7:0] a_146,
output reg [7:0] a_147,
output reg [7:0] a_148,
output reg [7:0] a_149,
output reg [7:0] a_150,
output reg [7:0] a_151,
output reg [7:0] a_152,
output reg [7:0] a_153,
output reg [7:0] a_154,
output reg [7:0] a_155,
output reg [7:0] a_156,
output reg [7:0] a_157,
output reg [7:0] a_158,
output reg [7:0] a_159,
output reg [7:0] a_160,
output reg [7:0] a_161,
output reg [7:0] a_162,
output reg [7:0] a_163,
output reg [7:0] a_164,
output reg [7:0] a_165,
output reg [7:0] a_166,
output reg [7:0] a_167,
output reg [7:0] a_168,
output reg [7:0] a_169,
output reg [7:0] a_170,
output reg [7:0] a_171,
output reg [7:0] a_172,
output reg [7:0] a_173,
output reg [7:0] a_174,
output reg [7:0] a_175,
output reg [7:0] a_176,
output reg [7:0] a_177,
output reg [7:0] a_178,
output reg [7:0] a_179,
output reg [7:0] a_180,
output reg [7:0] a_181,
output reg [7:0] a_182,
output reg [7:0] a_183,
output reg [7:0] a_184,
output reg [7:0] a_185,
output reg [7:0] a_186,
output reg [7:0] a_187,
output reg [7:0] a_188,
output reg [7:0] a_189,
output reg [7:0] a_190,
output reg [7:0] a_191,
output reg [7:0] a_192,
output reg [7:0] a_193,
output reg [7:0] a_194,
output reg [7:0] a_195,
output reg [7:0] a_196,
output reg [7:0] a_197,
output reg [7:0] a_198,
output reg [7:0] a_199,
output reg [7:0] a_200,
output reg [7:0] a_201,
output reg [7:0] a_202,
output reg [7:0] a_203,
output reg [7:0] a_204,
output reg [7:0] a_205,
output reg [7:0] a_206,
output reg [7:0] a_207,
output reg [7:0] a_208,
output reg [7:0] a_209,
output reg [7:0] a_210,
output reg [7:0] a_211,
output reg [7:0] a_212,
output reg [7:0] a_213,
output reg [7:0] a_214,
output reg [7:0] a_215,
output reg [7:0] a_216,
output reg [7:0] a_217,
output reg [7:0] a_218,
output reg [7:0] a_219,
output reg [7:0] a_220,
output reg [7:0] a_221,
output reg [7:0] a_222,
output reg [7:0] a_223,
output reg [7:0] a_224,
output reg [7:0] a_225,
output reg [7:0] a_226,
output reg [7:0] a_227,
output reg [7:0] a_228,
output reg [7:0] a_229,
output reg [7:0] a_230,
output reg [7:0] a_231,
output reg [7:0] a_232,
output reg [7:0] a_233,
output reg [7:0] a_234,
output reg [7:0] a_235,
output reg [7:0] a_236,
output reg [7:0] a_237,
output reg [7:0] a_238,
output reg [7:0] a_239,
output reg [7:0] a_240,
output reg [7:0] a_241,
output reg [7:0] a_242,
output reg [7:0] a_243,
output reg [7:0] a_244,
output reg [7:0] a_245,
output reg [7:0] a_246,
output reg [7:0] a_247,
output reg [7:0] a_248,
output reg [7:0] a_249,
output reg [7:0] a_250,
output reg [7:0] a_251,
output reg [7:0] a_252,
output reg [7:0] a_253,
output reg [7:0] a_254,
output reg [7:0] a_255,
output reg [7:0] a_256,
output reg [7:0] a_257,
output reg [7:0] a_258,
output reg [7:0] a_259,
output reg [7:0] a_260,
output reg [7:0] a_261,
output reg [7:0] a_262,
output reg [7:0] a_263,
output reg [7:0] a_264,
output reg [7:0] a_265,
output reg [7:0] a_266,
output reg [7:0] a_267,
output reg [7:0] a_268,
output reg [7:0] a_269,
output reg [7:0] a_270,
output reg [7:0] a_271,
output reg [7:0] a_272,
output reg [7:0] a_273,
output reg [7:0] a_274,
output reg [7:0] a_275,
output reg [7:0] a_276,
output reg [7:0] a_277,
output reg [7:0] a_278,
output reg [7:0] a_279,
output reg [7:0] a_280,
output reg [7:0] a_281,
output reg [7:0] a_282,
output reg [7:0] a_283,
output reg [7:0] a_284,
output reg [7:0] a_285,
output reg [7:0] a_286,
output reg [7:0] a_287,
output reg [7:0] a_288
);

reg [8:0] counter=0;
always @(posedge clk)
begin 
    case (counter)
    9'h00: a_1 <= a;
    9'h01: a_2 <= a;
    9'h02: a_3 <= a;
    9'h03: a_4 <= a;
    9'h04: a_5 <= a;
    9'h05: a_6 <= a;
    9'h06: a_7 <= a;
    9'h07: a_8 <= a;
    9'h08: a_9 <= a;
    9'h09: a_10 <= a;
    9'h0A: a_11 <= a;
    9'h0B: a_12 <= a;
    9'h0C: a_13 <= a;
    9'h0D: a_14 <= a;
    9'h0E: a_15 <= a;
    9'h0F: a_16 <= a;
    9'h10: a_17 <= a;
    9'h11: a_18 <= a;
    9'h12: a_19 <= a;
    9'h13: a_20 <= a;
    9'h14: a_21 <= a;
    9'h15: a_22 <= a;
    9'h16: a_23 <= a;
    9'h17: a_24 <= a;
    9'h18: a_25 <= a;
    9'h19: a_26 <= a;
    9'h1A: a_27 <= a;
    9'h1B: a_28 <= a;
    9'h1C: a_29 <= a;
    9'h1D: a_30 <= a;
    9'h1E: a_31 <= a;
    9'h1F: a_32 <= a;
    9'h20: a_33 <= a;
    9'h21: a_34 <= a;
    9'h22: a_35 <= a;
    9'h23: a_36 <= a;
    9'h24: a_37 <= a;
    9'h25: a_38 <= a;
    9'h26: a_39 <= a;
    9'h27: a_40 <= a;
    9'h28: a_41 <= a;
    9'h29: a_42 <= a;
    9'h2A: a_43 <= a;
    9'h2B: a_44 <= a;
    9'h2C: a_45 <= a;
    9'h2D: a_46 <= a;
    9'h2E: a_47 <= a;
    9'h2F: a_48 <= a;
    9'h30: a_49 <= a;
    9'h31: a_50 <= a;
    9'h32: a_51 <= a;
    9'h33: a_52 <= a;
    9'h34: a_53 <= a;
    9'h35: a_54 <= a;
    9'h36: a_55 <= a;
    9'h37: a_56 <= a;
    9'h38: a_57 <= a;
    9'h39: a_58 <= a;
    9'h3A: a_59 <= a;
    9'h3B: a_60 <= a;
    9'h3C: a_61 <= a;
    9'h3D: a_62 <= a;
    9'h3E: a_63 <= a;
    9'h3F: a_64 <= a;
    9'h40: a_65 <= a;
    9'h41: a_66 <= a;
    9'h42: a_67 <= a;
    9'h43: a_68 <= a;
    9'h44: a_69 <= a;
    9'h45: a_70 <= a;
    9'h46: a_71 <= a;
    9'h47: a_72 <= a;
    9'h48: a_73 <= a;
    9'h49: a_74 <= a;
    9'h4A: a_75 <= a;
    9'h4B: a_76 <= a;
    9'h4C: a_77 <= a;
    9'h4D: a_78 <= a;
    9'h4E: a_79 <= a;
    9'h4F: a_80 <= a;
    9'h50: a_81 <= a;
    9'h51: a_82 <= a;
    9'h52: a_83 <= a;
    9'h53: a_84 <= a;
    9'h54: a_85 <= a;
    9'h55: a_86 <= a;
    9'h56: a_87 <= a;
    9'h57: a_88 <= a;
    9'h58: a_89 <= a;
    9'h59: a_90 <= a;
    9'h5A: a_91 <= a;
    9'h5B: a_92 <= a;
    9'h5C: a_93 <= a;
    9'h5D: a_94 <= a;
    9'h5E: a_95 <= a;
    9'h5F: a_96 <= a;
    9'h60: a_97 <= a;
    9'h61: a_98 <= a;
    9'h62: a_99 <= a;
    9'h63: a_100 <= a;
    9'h64: a_101 <= a;
    9'h65: a_102 <= a;
    9'h66: a_103 <= a;
    9'h67: a_104 <= a;
    9'h68: a_105 <= a;
    9'h69: a_106 <= a;
    9'h6A: a_107 <= a;
    9'h6B: a_108 <= a;
    9'h6C: a_109 <= a;
    9'h6D: a_110 <= a;
    9'h6E: a_111 <= a;
    9'h6F: a_112 <= a;
    9'h70: a_113 <= a;
    9'h71: a_114 <= a;
    9'h72: a_115 <= a;
    9'h73: a_116 <= a;
    9'h74: a_117 <= a;
    9'h75: a_118 <= a;
    9'h76: a_119 <= a;
    9'h77: a_120 <= a;
    9'h78: a_121 <= a;
    9'h79: a_122 <= a;
    9'h7A: a_123 <= a;
    9'h7B: a_124 <= a;
    9'h7C: a_125 <= a;
    9'h7D: a_126 <= a;
    9'h7E: a_127 <= a;
    9'h7F: a_128 <= a;
    9'h80: a_129 <= a;
    9'h81: a_130 <= a;
    9'h82: a_131 <= a;
    9'h83: a_132 <= a;
    9'h84: a_133 <= a;
    9'h85: a_134 <= a;
    9'h86: a_135 <= a;
    9'h87: a_136 <= a;
    9'h88: a_137 <= a;
    9'h89: a_138 <= a;
    9'h8A: a_139 <= a;
    9'h8B: a_140 <= a;
    9'h8C: a_141 <= a;
    9'h8D: a_142 <= a;
    9'h8E: a_143 <= a;
    9'h8F: a_144 <= a;
    9'h90: a_145 <= a;
    9'h91: a_146 <= a;
    9'h92: a_147 <= a;
    9'h93: a_148 <= a;
    9'h94: a_149 <= a;
    9'h95: a_150 <= a;
    9'h96: a_151 <= a;
    9'h97: a_152 <= a;
    9'h98: a_153 <= a;
    9'h99: a_154 <= a;
    9'h9A: a_155 <= a;
    9'h9B: a_156 <= a;
    9'h9C: a_157 <= a;
    9'h9D: a_158 <= a;
    9'h9E: a_159 <= a;
    9'h9F: a_160 <= a;
    9'hA0: a_161 <= a;
    9'hA1: a_162 <= a;
    9'hA2: a_163 <= a;
    9'hA3: a_164 <= a;
    9'hA4: a_165 <= a;
    9'hA5: a_166 <= a;
    9'hA6: a_167 <= a;
    9'hA7: a_168 <= a;
    9'hA8: a_169 <= a;
    9'hA9: a_170 <= a;
    9'hAA: a_171 <= a;
    9'hAB: a_172 <= a;
    9'hAC: a_173 <= a;
    9'hAD: a_174 <= a;
    9'hAE: a_175 <= a;
    9'hAF: a_176 <= a;
    9'hB0: a_177 <= a;
    9'hB1: a_178 <= a;
    9'hB2: a_179 <= a;
    9'hB3: a_180 <= a;
    9'hB4: a_181 <= a;
    9'hB5: a_182 <= a;
    9'hB6: a_183 <= a;
    9'hB7: a_184 <= a;
    9'hB8: a_185 <= a;
    9'hB9: a_186 <= a;
    9'hBA: a_187 <= a;
    9'hBB: a_188 <= a;
    9'hBC: a_189 <= a;
    9'hBD: a_190 <= a;
    9'hBE: a_191 <= a;
    9'hBF: a_192 <= a;
    9'hC0: a_193 <= a;
    9'hC1: a_194 <= a;
    9'hC2: a_195 <= a;
    9'hC3: a_196 <= a;
    9'hC4: a_197 <= a;
    9'hC5: a_198 <= a;
    9'hC6: a_199 <= a;
    9'hC7: a_200 <= a;
    9'hC8: a_201 <= a;
    9'hC9: a_202 <= a;
    9'hCA: a_203 <= a;
    9'hCB: a_204 <= a;
    9'hCC: a_205 <= a;
    9'hCD: a_206 <= a;
    9'hCE: a_207 <= a;
    9'hCF: a_208 <= a;
    9'hD0: a_209 <= a;
    9'hD1: a_210 <= a;
    9'hD2: a_211 <= a;
    9'hD3: a_212 <= a;
    9'hD4: a_213 <= a;
    9'hD5: a_214 <= a;
    9'hD6: a_215 <= a;
    9'hD7: a_216 <= a;
    9'hD8: a_217 <= a;
    9'hD9: a_218 <= a;
    9'hDA: a_219 <= a;
    9'hDB: a_220 <= a;
    9'hDC: a_221 <= a;
    9'hDD: a_222 <= a;
    9'hDE: a_223 <= a;
    9'hDF: a_224 <= a;
    9'hE0: a_225 <= a;
    9'hE1: a_226 <= a;
    9'hE2: a_227 <= a;
    9'hE3: a_228 <= a;
    9'hE4: a_229 <= a;
    9'hE5: a_230 <= a;
    9'hE6: a_231 <= a;
    9'hE7: a_232 <= a;
    9'hE8: a_233 <= a;
    9'hE9: a_234 <= a;
    9'hEA: a_235 <= a;
    9'hEB: a_236 <= a;
    9'hEC: a_237 <= a;
    9'hED: a_238 <= a;
    9'hEE: a_239 <= a;
    9'hEF: a_240 <= a;
    9'hF0: a_241 <= a;
    9'hF1: a_242 <= a;
    9'hF2: a_243 <= a;
    9'hF3: a_244 <= a;
    9'hF4: a_245 <= a;
    9'hF5: a_246 <= a;
    9'hF6: a_247 <= a;
    9'hF7: a_248 <= a;
    9'hF8: a_249 <= a;
    9'hF9: a_250 <= a;
    9'hFA: a_251 <= a;
    9'hFB: a_252 <= a;
    9'hFC: a_253 <= a;
    9'hFD: a_254 <= a;
    9'hFE: a_255 <= a;
    9'hFF: a_256 <= a;
    9'h100: a_257 <= a;
    9'h101: a_258 <= a;
    9'h102: a_259 <= a;
    9'h103: a_260 <= a;
    9'h104: a_261 <= a;
    9'h105: a_262 <= a;
    9'h106: a_263 <= a;
    9'h107: a_264 <= a;
    9'h108: a_265 <= a;
    9'h109: a_266 <= a;
    9'h10A: a_267 <= a;
    9'h10B: a_268 <= a;
    9'h10C: a_269 <= a;
    9'h10D: a_270 <= a;
    9'h10E: a_271 <= a;
    9'h10F: a_272 <= a;
    9'h110: a_273 <= a;
    9'h111: a_274 <= a;
    9'h112: a_275 <= a;
    9'h113: a_276 <= a;
    9'h114: a_277 <= a;
    9'h115: a_278 <= a;
    9'h116: a_279 <= a;
    9'h117: a_280 <= a;
    9'h118: a_281 <= a;
    9'h119: a_282 <= a;
    9'h11A: a_283 <= a;
    9'h11B: a_284 <= a;
    9'h11C: a_285 <= a;
    9'h11D: a_286 <= a;
    9'h11E: a_287 <= a;
    9'h11F: a_288 <= a;
    default:a_1<=a;
endcase

   counter<=counter+1;
   end
   
   endmodule

    
