`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.10.2023 14:44:30
// Design Name: 
// Module Name: fa
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fa(
input A,
input B,
input Cin,
output Cout,
output Y
    );

wire [1:0] temp;
assign temp=A+B+Cin;
assign Y=temp[0];
assign Cout=temp[1];


//  assign Y=A^B^Cin;
//  assign Cout=(A^B)&Cin | A&B;
endmodule
